///Calculating Leftmost Set bit//////////////////
Approach-1: Right Shift the Number till its greater than 0 (>0) . 
